-- QSYS_SC_TEI0026.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity QSYS_SC_TEI0026 is
	port (
		clk_in_clk              : in  std_logic                    := '0';             --           clk_in.clk
		pio_in_dip_sw_export    : in  std_logic_vector(3 downto 0) := (others => '0'); --    pio_in_dip_sw.export
		pio_in_usr_export       : in  std_logic_vector(2 downto 0) := (others => '0'); --       pio_in_usr.export
		pio_out_user_led_export : out std_logic_vector(3 downto 0);                    -- pio_out_user_led.export
		pio_out_vdd1_export     : out std_logic_vector(4 downto 0);                    --     pio_out_vdd1.export
		pio_out_vdd2_export     : out std_logic_vector(5 downto 0);                    --     pio_out_vdd2.export
		pio_out_vdd3_export     : out std_logic_vector(4 downto 0);                    --     pio_out_vdd3.export
		reset_reset_n           : in  std_logic                    := '0';             --            reset.reset_n
		uart_rxd                : in  std_logic                    := '0';             --             uart.rxd
		uart_txd                : out std_logic                                        --                 .txd
	);
end entity QSYS_SC_TEI0026;

architecture rtl of QSYS_SC_TEI0026 is
	component QSYS_SC_TEI0026_nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component QSYS_SC_TEI0026_nios2;

	component QSYS_SC_TEI0026_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component QSYS_SC_TEI0026_onchip_ram;

	component QSYS_SC_TEI0026_pio_in_dip_sw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component QSYS_SC_TEI0026_pio_in_dip_sw;

	component QSYS_SC_TEI0026_pio_in_usr is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component QSYS_SC_TEI0026_pio_in_usr;

	component QSYS_SC_TEI0026_pio_out_user_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component QSYS_SC_TEI0026_pio_out_user_led;

	component QSYS_SC_TEI0026_pio_out_vdd1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(4 downto 0)                      -- export
		);
	end component QSYS_SC_TEI0026_pio_out_vdd1;

	component QSYS_SC_TEI0026_pio_out_vdd2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component QSYS_SC_TEI0026_pio_out_vdd2;

	component QSYS_SC_TEI0026_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component QSYS_SC_TEI0026_pll;

	component QSYS_SC_TEI0026_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component QSYS_SC_TEI0026_uart;

	component QSYS_SC_TEI0026_mm_interconnect_0 is
		port (
			clk_in_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			nios2_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_data_master_address                             : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                                : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_write                               : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address                      : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_debug_mem_slave_address                         : out std_logic_vector(8 downto 0);                     -- address
			nios2_debug_mem_slave_write                           : out std_logic;                                        -- write
			nios2_debug_mem_slave_read                            : out std_logic;                                        -- read
			nios2_debug_mem_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_debug_mem_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_debug_mem_slave_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_debug_mem_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			nios2_debug_mem_slave_debugaccess                     : out std_logic;                                        -- debugaccess
			onchip_ram_s1_address                                 : out std_logic_vector(12 downto 0);                    -- address
			onchip_ram_s1_write                                   : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                   : out std_logic;                                        -- clken
			pio_in_dip_sw_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			pio_in_dip_sw_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_in_usr_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_in_usr_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_user_led_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			pio_out_user_led_s1_write                             : out std_logic;                                        -- write
			pio_out_user_led_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_user_led_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_user_led_s1_chipselect                        : out std_logic;                                        -- chipselect
			pio_out_vdd1_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pio_out_vdd1_s1_write                                 : out std_logic;                                        -- write
			pio_out_vdd1_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_vdd1_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_vdd1_s1_chipselect                            : out std_logic;                                        -- chipselect
			pio_out_vdd2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pio_out_vdd2_s1_write                                 : out std_logic;                                        -- write
			pio_out_vdd2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_vdd2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_vdd2_s1_chipselect                            : out std_logic;                                        -- chipselect
			pio_out_vdd3_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pio_out_vdd3_s1_write                                 : out std_logic;                                        -- write
			pio_out_vdd3_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_vdd3_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_vdd3_s1_chipselect                            : out std_logic;                                        -- chipselect
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			uart_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                                         : out std_logic;                                        -- write
			uart_s1_read                                          : out std_logic;                                        -- read
			uart_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                                 : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component QSYS_SC_TEI0026_mm_interconnect_0;

	component QSYS_SC_TEI0026_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component QSYS_SC_TEI0026_irq_mapper;

	component qsys_sc_tei0026_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsys_sc_tei0026_rst_controller;

	component qsys_sc_tei0026_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsys_sc_tei0026_rst_controller_001;

	signal pll_c0_clk                                            : std_logic;                     -- pll:c0 -> [irq_mapper:clk, mm_interconnect_0:pll_c0_clk, nios2:clk, onchip_ram:clk, pio_in_dip_sw:clk, pio_in_usr:clk, pio_out_user_led:clk, pio_out_vdd1:clk, pio_out_vdd2:clk, pio_out_vdd3:clk, rst_controller:clk, uart:clk]
	signal nios2_data_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                         : std_logic;                     -- nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_address                             : std_logic_vector(16 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_byteenable                          : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal nios2_data_master_read                                : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_write                               : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_writedata                           : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal nios2_instruction_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                  : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                      : std_logic_vector(16 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                         : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal mm_interconnect_0_nios2_debug_mem_slave_readdata      : std_logic_vector(31 downto 0); -- nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_debug_mem_slave_waitrequest   : std_logic;                     -- nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_debug_mem_slave_debugaccess   : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_debug_mem_slave_address       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_debug_mem_slave_read          : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_debug_mem_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_debug_mem_slave_write         : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_debug_mem_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata              : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                  : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                 : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect            : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata              : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address               : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                 : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                 : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_uart_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                    : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                        : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer               : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                       : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal mm_interconnect_0_pio_in_usr_s1_readdata              : std_logic_vector(31 downto 0); -- pio_in_usr:readdata -> mm_interconnect_0:pio_in_usr_s1_readdata
	signal mm_interconnect_0_pio_in_usr_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_in_usr_s1_address -> pio_in_usr:address
	signal mm_interconnect_0_pio_in_dip_sw_s1_readdata           : std_logic_vector(31 downto 0); -- pio_in_dip_sw:readdata -> mm_interconnect_0:pio_in_dip_sw_s1_readdata
	signal mm_interconnect_0_pio_in_dip_sw_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_in_dip_sw_s1_address -> pio_in_dip_sw:address
	signal mm_interconnect_0_pio_out_vdd1_s1_chipselect          : std_logic;                     -- mm_interconnect_0:pio_out_vdd1_s1_chipselect -> pio_out_vdd1:chipselect
	signal mm_interconnect_0_pio_out_vdd1_s1_readdata            : std_logic_vector(31 downto 0); -- pio_out_vdd1:readdata -> mm_interconnect_0:pio_out_vdd1_s1_readdata
	signal mm_interconnect_0_pio_out_vdd1_s1_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_vdd1_s1_address -> pio_out_vdd1:address
	signal mm_interconnect_0_pio_out_vdd1_s1_write               : std_logic;                     -- mm_interconnect_0:pio_out_vdd1_s1_write -> mm_interconnect_0_pio_out_vdd1_s1_write:in
	signal mm_interconnect_0_pio_out_vdd1_s1_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_vdd1_s1_writedata -> pio_out_vdd1:writedata
	signal mm_interconnect_0_pio_out_vdd2_s1_chipselect          : std_logic;                     -- mm_interconnect_0:pio_out_vdd2_s1_chipselect -> pio_out_vdd2:chipselect
	signal mm_interconnect_0_pio_out_vdd2_s1_readdata            : std_logic_vector(31 downto 0); -- pio_out_vdd2:readdata -> mm_interconnect_0:pio_out_vdd2_s1_readdata
	signal mm_interconnect_0_pio_out_vdd2_s1_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_vdd2_s1_address -> pio_out_vdd2:address
	signal mm_interconnect_0_pio_out_vdd2_s1_write               : std_logic;                     -- mm_interconnect_0:pio_out_vdd2_s1_write -> mm_interconnect_0_pio_out_vdd2_s1_write:in
	signal mm_interconnect_0_pio_out_vdd2_s1_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_vdd2_s1_writedata -> pio_out_vdd2:writedata
	signal mm_interconnect_0_pio_out_vdd3_s1_chipselect          : std_logic;                     -- mm_interconnect_0:pio_out_vdd3_s1_chipselect -> pio_out_vdd3:chipselect
	signal mm_interconnect_0_pio_out_vdd3_s1_readdata            : std_logic_vector(31 downto 0); -- pio_out_vdd3:readdata -> mm_interconnect_0:pio_out_vdd3_s1_readdata
	signal mm_interconnect_0_pio_out_vdd3_s1_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_vdd3_s1_address -> pio_out_vdd3:address
	signal mm_interconnect_0_pio_out_vdd3_s1_write               : std_logic;                     -- mm_interconnect_0:pio_out_vdd3_s1_write -> mm_interconnect_0_pio_out_vdd3_s1_write:in
	signal mm_interconnect_0_pio_out_vdd3_s1_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_vdd3_s1_writedata -> pio_out_vdd3:writedata
	signal mm_interconnect_0_pio_out_user_led_s1_chipselect      : std_logic;                     -- mm_interconnect_0:pio_out_user_led_s1_chipselect -> pio_out_user_led:chipselect
	signal mm_interconnect_0_pio_out_user_led_s1_readdata        : std_logic_vector(31 downto 0); -- pio_out_user_led:readdata -> mm_interconnect_0:pio_out_user_led_s1_readdata
	signal mm_interconnect_0_pio_out_user_led_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_user_led_s1_address -> pio_out_user_led:address
	signal mm_interconnect_0_pio_out_user_led_s1_write           : std_logic;                     -- mm_interconnect_0:pio_out_user_led_s1_write -> mm_interconnect_0_pio_out_user_led_s1_write:in
	signal mm_interconnect_0_pio_out_user_led_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_user_led_s1_writedata -> pio_out_user_led:writedata
	signal irq_mapper_receiver0_irq                              : std_logic;                     -- uart:irq -> irq_mapper:receiver0_irq
	signal nios2_irq_irq                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:irq
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                    : std_logic;                     -- rst_controller:reset_req -> [nios2:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal nios2_debug_reset_request_reset                       : std_logic;                     -- nios2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                    : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                               : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_uart_s1_read_ports_inv              : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal mm_interconnect_0_pio_out_vdd1_s1_write_ports_inv     : std_logic;                     -- mm_interconnect_0_pio_out_vdd1_s1_write:inv -> pio_out_vdd1:write_n
	signal mm_interconnect_0_pio_out_vdd2_s1_write_ports_inv     : std_logic;                     -- mm_interconnect_0_pio_out_vdd2_s1_write:inv -> pio_out_vdd2:write_n
	signal mm_interconnect_0_pio_out_vdd3_s1_write_ports_inv     : std_logic;                     -- mm_interconnect_0_pio_out_vdd3_s1_write:inv -> pio_out_vdd3:write_n
	signal mm_interconnect_0_pio_out_user_led_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_pio_out_user_led_s1_write:inv -> pio_out_user_led:write_n
	signal rst_controller_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [nios2:reset_n, pio_in_dip_sw:reset_n, pio_in_usr:reset_n, pio_out_user_led:reset_n, pio_out_vdd1:reset_n, pio_out_vdd2:reset_n, pio_out_vdd3:reset_n, uart:reset_n]

begin

	nios2 : component QSYS_SC_TEI0026_nios2
		port map (
			clk                                 => pll_c0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	onchip_ram : component QSYS_SC_TEI0026_onchip_ram
		port map (
			clk        => pll_c0_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pio_in_dip_sw : component QSYS_SC_TEI0026_pio_in_dip_sw
		port map (
			clk      => pll_c0_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_pio_in_dip_sw_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_in_dip_sw_s1_readdata, --                    .readdata
			in_port  => pio_in_dip_sw_export                         -- external_connection.export
		);

	pio_in_usr : component QSYS_SC_TEI0026_pio_in_usr
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pio_in_usr_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_in_usr_s1_readdata, --                    .readdata
			in_port  => pio_in_usr_export                         -- external_connection.export
		);

	pio_out_user_led : component QSYS_SC_TEI0026_pio_out_user_led
		port map (
			clk        => pll_c0_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_pio_out_user_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_user_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_user_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_user_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_user_led_s1_readdata,        --                    .readdata
			out_port   => pio_out_user_led_export                                -- external_connection.export
		);

	pio_out_vdd1 : component QSYS_SC_TEI0026_pio_out_vdd1
		port map (
			clk        => pll_c0_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_pio_out_vdd1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_vdd1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_vdd1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_vdd1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_vdd1_s1_readdata,        --                    .readdata
			out_port   => pio_out_vdd1_export                                -- external_connection.export
		);

	pio_out_vdd2 : component QSYS_SC_TEI0026_pio_out_vdd2
		port map (
			clk        => pll_c0_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_pio_out_vdd2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_vdd2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_vdd2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_vdd2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_vdd2_s1_readdata,        --                    .readdata
			out_port   => pio_out_vdd2_export                                -- external_connection.export
		);

	pio_out_vdd3 : component QSYS_SC_TEI0026_pio_out_vdd1
		port map (
			clk        => pll_c0_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_pio_out_vdd3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_vdd3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_vdd3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_vdd3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_vdd3_s1_readdata,        --                    .readdata
			out_port   => pio_out_vdd3_export                                -- external_connection.export
		);

	pll : component QSYS_SC_TEI0026_pll
		port map (
			clk                => clk_in_clk,                                --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c1                 => open,                                      --           (terminated)
			c2                 => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	uart : component QSYS_SC_TEI0026_uart
		port map (
			clk           => pll_c0_clk,                                --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => uart_rxd,                                  -- external_connection.export
			txd           => uart_txd,                                  --                    .export
			irq           => irq_mapper_receiver0_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component QSYS_SC_TEI0026_mm_interconnect_0
		port map (
			clk_in_clk_clk                                        => clk_in_clk,                                          --                                      clk_in_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                          --                                          pll_c0.clk
			nios2_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                      --               nios2_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                  -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_data_master_address                             => nios2_data_master_address,                           --                               nios2_data_master.address
			nios2_data_master_waitrequest                         => nios2_data_master_waitrequest,                       --                                                .waitrequest
			nios2_data_master_byteenable                          => nios2_data_master_byteenable,                        --                                                .byteenable
			nios2_data_master_read                                => nios2_data_master_read,                              --                                                .read
			nios2_data_master_readdata                            => nios2_data_master_readdata,                          --                                                .readdata
			nios2_data_master_write                               => nios2_data_master_write,                             --                                                .write
			nios2_data_master_writedata                           => nios2_data_master_writedata,                         --                                                .writedata
			nios2_data_master_debugaccess                         => nios2_data_master_debugaccess,                       --                                                .debugaccess
			nios2_instruction_master_address                      => nios2_instruction_master_address,                    --                        nios2_instruction_master.address
			nios2_instruction_master_waitrequest                  => nios2_instruction_master_waitrequest,                --                                                .waitrequest
			nios2_instruction_master_read                         => nios2_instruction_master_read,                       --                                                .read
			nios2_instruction_master_readdata                     => nios2_instruction_master_readdata,                   --                                                .readdata
			nios2_debug_mem_slave_address                         => mm_interconnect_0_nios2_debug_mem_slave_address,     --                           nios2_debug_mem_slave.address
			nios2_debug_mem_slave_write                           => mm_interconnect_0_nios2_debug_mem_slave_write,       --                                                .write
			nios2_debug_mem_slave_read                            => mm_interconnect_0_nios2_debug_mem_slave_read,        --                                                .read
			nios2_debug_mem_slave_readdata                        => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                                                .readdata
			nios2_debug_mem_slave_writedata                       => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                                                .writedata
			nios2_debug_mem_slave_byteenable                      => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                                                .byteenable
			nios2_debug_mem_slave_waitrequest                     => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                                                .waitrequest
			nios2_debug_mem_slave_debugaccess                     => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                                                .debugaccess
			onchip_ram_s1_address                                 => mm_interconnect_0_onchip_ram_s1_address,             --                                   onchip_ram_s1.address
			onchip_ram_s1_write                                   => mm_interconnect_0_onchip_ram_s1_write,               --                                                .write
			onchip_ram_s1_readdata                                => mm_interconnect_0_onchip_ram_s1_readdata,            --                                                .readdata
			onchip_ram_s1_writedata                               => mm_interconnect_0_onchip_ram_s1_writedata,           --                                                .writedata
			onchip_ram_s1_byteenable                              => mm_interconnect_0_onchip_ram_s1_byteenable,          --                                                .byteenable
			onchip_ram_s1_chipselect                              => mm_interconnect_0_onchip_ram_s1_chipselect,          --                                                .chipselect
			onchip_ram_s1_clken                                   => mm_interconnect_0_onchip_ram_s1_clken,               --                                                .clken
			pio_in_dip_sw_s1_address                              => mm_interconnect_0_pio_in_dip_sw_s1_address,          --                                pio_in_dip_sw_s1.address
			pio_in_dip_sw_s1_readdata                             => mm_interconnect_0_pio_in_dip_sw_s1_readdata,         --                                                .readdata
			pio_in_usr_s1_address                                 => mm_interconnect_0_pio_in_usr_s1_address,             --                                   pio_in_usr_s1.address
			pio_in_usr_s1_readdata                                => mm_interconnect_0_pio_in_usr_s1_readdata,            --                                                .readdata
			pio_out_user_led_s1_address                           => mm_interconnect_0_pio_out_user_led_s1_address,       --                             pio_out_user_led_s1.address
			pio_out_user_led_s1_write                             => mm_interconnect_0_pio_out_user_led_s1_write,         --                                                .write
			pio_out_user_led_s1_readdata                          => mm_interconnect_0_pio_out_user_led_s1_readdata,      --                                                .readdata
			pio_out_user_led_s1_writedata                         => mm_interconnect_0_pio_out_user_led_s1_writedata,     --                                                .writedata
			pio_out_user_led_s1_chipselect                        => mm_interconnect_0_pio_out_user_led_s1_chipselect,    --                                                .chipselect
			pio_out_vdd1_s1_address                               => mm_interconnect_0_pio_out_vdd1_s1_address,           --                                 pio_out_vdd1_s1.address
			pio_out_vdd1_s1_write                                 => mm_interconnect_0_pio_out_vdd1_s1_write,             --                                                .write
			pio_out_vdd1_s1_readdata                              => mm_interconnect_0_pio_out_vdd1_s1_readdata,          --                                                .readdata
			pio_out_vdd1_s1_writedata                             => mm_interconnect_0_pio_out_vdd1_s1_writedata,         --                                                .writedata
			pio_out_vdd1_s1_chipselect                            => mm_interconnect_0_pio_out_vdd1_s1_chipselect,        --                                                .chipselect
			pio_out_vdd2_s1_address                               => mm_interconnect_0_pio_out_vdd2_s1_address,           --                                 pio_out_vdd2_s1.address
			pio_out_vdd2_s1_write                                 => mm_interconnect_0_pio_out_vdd2_s1_write,             --                                                .write
			pio_out_vdd2_s1_readdata                              => mm_interconnect_0_pio_out_vdd2_s1_readdata,          --                                                .readdata
			pio_out_vdd2_s1_writedata                             => mm_interconnect_0_pio_out_vdd2_s1_writedata,         --                                                .writedata
			pio_out_vdd2_s1_chipselect                            => mm_interconnect_0_pio_out_vdd2_s1_chipselect,        --                                                .chipselect
			pio_out_vdd3_s1_address                               => mm_interconnect_0_pio_out_vdd3_s1_address,           --                                 pio_out_vdd3_s1.address
			pio_out_vdd3_s1_write                                 => mm_interconnect_0_pio_out_vdd3_s1_write,             --                                                .write
			pio_out_vdd3_s1_readdata                              => mm_interconnect_0_pio_out_vdd3_s1_readdata,          --                                                .readdata
			pio_out_vdd3_s1_writedata                             => mm_interconnect_0_pio_out_vdd3_s1_writedata,         --                                                .writedata
			pio_out_vdd3_s1_chipselect                            => mm_interconnect_0_pio_out_vdd3_s1_chipselect,        --                                                .chipselect
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,             --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,               --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,            --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,           --                                                .writedata
			uart_s1_address                                       => mm_interconnect_0_uart_s1_address,                   --                                         uart_s1.address
			uart_s1_write                                         => mm_interconnect_0_uart_s1_write,                     --                                                .write
			uart_s1_read                                          => mm_interconnect_0_uart_s1_read,                      --                                                .read
			uart_s1_readdata                                      => mm_interconnect_0_uart_s1_readdata,                  --                                                .readdata
			uart_s1_writedata                                     => mm_interconnect_0_uart_s1_writedata,                 --                                                .writedata
			uart_s1_begintransfer                                 => mm_interconnect_0_uart_s1_begintransfer,             --                                                .begintransfer
			uart_s1_chipselect                                    => mm_interconnect_0_uart_s1_chipselect                 --                                                .chipselect
		);

	irq_mapper : component QSYS_SC_TEI0026_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_irq_irq                   --    sender.irq
		);

	rst_controller : component qsys_sc_tei0026_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component qsys_sc_tei0026_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => clk_in_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	mm_interconnect_0_pio_out_vdd1_s1_write_ports_inv <= not mm_interconnect_0_pio_out_vdd1_s1_write;

	mm_interconnect_0_pio_out_vdd2_s1_write_ports_inv <= not mm_interconnect_0_pio_out_vdd2_s1_write;

	mm_interconnect_0_pio_out_vdd3_s1_write_ports_inv <= not mm_interconnect_0_pio_out_vdd3_s1_write;

	mm_interconnect_0_pio_out_user_led_s1_write_ports_inv <= not mm_interconnect_0_pio_out_user_led_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of QSYS_SC_TEI0026
